/*
Author: Prerak Chaudhari
Student Number: 1005114760

Date: September 26th, 2019
*/

module lab2part1(SW, LEDR);
	input [9:0] SW;
	output [9:0] LEDR;
	
	assign LEDR = SW;
endmodule